Simulation of the symmetrical OTA designed with the sEKV model by C. Enz

.include ekv018va.par ; model file for EKV2.6
.include size_bias.par ; Size and bias values
.include Symmetrical_OTA.net ; Circuit netlist

.control
 op
 save inoise_spectrum onoise_spectrum
 + onoise_n1a onoise_n1b onoise_n1a_thermal onoise_n1b_thermal onoise_n1a_flicker onoise_n1b_flicker
 + onoise_n2a onoise_n2b onoise_n2c onoise_n2d onoise_n2a_thermal onoise_n2b_thermal onoise_n2c_thermal onoise_n2d_thermal onoise_n2a_flicker onoise_n2b_flicker onoise_n2c_flicker onoise_n2d_flicker
 + onoise_n3a onoise_n3b onoise_n3a_thermal onoise_n3b_thermal onoise_n3a_flicker onoise_n3b_flicker
 + onoise_n4 onoise_n4_thermal onoise_n4_flicker
 + onoise_n7 onoise_n7_thermal onoise_n7_flicker
 noise V(out) Vid dec 41 1 100MEG 1
 setplot noise1
 write $inputdir/Symmetrical_OTA.nz.raw
 set wr_singlescale
 set wr_vecnames
 wrdata $inputdir/Symmetrical_OTA.nz.dat inoise_spectrum onoise_spectrum
.endc
.end
