Simulation of the CS stage optimized for GBW and DC gain

.include ekv018va.par ; model file for EKV2.6
.include size_bias.par ; Size and bias values
.include CS_GBW_Adc.net ; Circuit netlist

.control
 save @N1[Id] @N1[Ispec] @N1[IC] @N1[n0] @N1[gm] @N1[gms] @N1[gds] @N1[gmbs] @N1[Rn] @N1[Vnth] @N1[gamman] @N1[Vnfl] @N1[Vdsat]
 save @N2[Id] @N2[Ispec] @N2[IC] @N2[n0] @N2[gm] @N2[gms] @N2[gds] @N2[gmbs] @N2[Rn] @N2[Vnth] @N2[gamman] @N2[Vnfl] @N2[Vdsat]
 op
 wrnodev $inputdir/CS_GBW_Adc.op.ic
 set wr_singlescale
 set wr_vecnames
 wrdata $inputdir/CS_GBW_Adc.op.dat @N1[Id] @N1[Ispec] @N1[IC] @N1[Vdsat] @N1[n0] @N1[gm] @N1[gms] @N1[gds] @N1[gmbs] @N1[Rn] @N1[Vnth] @N1[gamman] @N1[Vnfl]
 set appendwrite
 wrdata $inputdir/CS_GBW_Adc.op.dat @N2[Id] @N2[Ispec] @N2[IC] @N2[Vdsat] @N2[n0] @N2[gm] @N2[gms] @N2[gds] @N2[gmbs] @N2[Rn] @N2[Vnth] @N2[gamman] @N2[Vnfl]
.endc
.end
