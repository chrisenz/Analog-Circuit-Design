Simulation of the symmetrical OTA designed with the EKV 2.6 model

.include ekv018va.par ; model file for EKV2.6
.include size_bias.par ; Size and bias values
.include Miller_OTA.net ; Circuit netlist

.control
 op
 save v(out)
 write $inputdir/Miller_OTA.ac.op
* reset all
 ac dec 41 100m 100MEG
 let AmagdB=vdb(out)
 let Aphdeg=180/PI*vp(out)
 meas ac Adc max AmagdB
 meas ac GBW when AmagdB=0
 meas ac PGBW find Aphdeg at=GBW
 set wr_singlescale
 set wr_vecnames
 wrdata $inputdir/Miller_OTA.ac.dat AmagdB Aphdeg
.endc
.end
